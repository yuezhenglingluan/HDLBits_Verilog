module top_module(
    input clk,
    input load,
    input [511:0] data,
    output [511:0] q ); 

endmodule
